
module control(input [2:0] opcode, 
output reg jump, branch, memwrite, regwrite
 );
 

