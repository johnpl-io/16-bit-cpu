module controller()

reg [15:0] instruction
reg [15:0] a