module controller()

reg [15:0] instruction;
reg [15:0] A, B;
reg [2:0] ALU_Code;